
.PARAM VDD = 1 VGS = 1 LN = 0.05U LP = 0.05U WN = 1U WP = 0.5U
M1 VOUT VIN 0 0 N_50n L = LN W = WN
M2 VOUT VIN VDD VDD P_50n L = LP W = WP
.INCLUDE 'C:\sdsy\model1\rf018.l'

VDD VDD 0 VDD
VIN VIN 0 VGS

.DC VIN 0 1 0.001

.PRINT v(VIN) v(VOUT)

.OPTION LIST NODE BRIEF=1 
.OPTION POST=3

.ALTER
.PARAM WN = 1.5U
.ALTER
.PARAM WN = 1U WP = 1U


.END