* .PARAM VDD = 1 VGS = 1 LN = 0.05U LP = 0.05U WN = 1U WP = 0.5U
* M1 VOUT VIN 0 0 N_50n L = LN W = WN
* M2 VOUT VIN VDD VDD P_50n L = LP W = WP
* C1 
.PARAM VDD = 1.8
M1 V1 VIN VDD VDD PCH L = 0.18U W = 15U
V1 V1 0 1.6
VIN VIN 0 1.8

VDD VDD 0 VDD
.DC VIN 0 1.8 0.001
.PRINT M1_VTH = par('lv9(M1)')

.OPTION LIST NODE BRIEF=1 
.OPTION POST=3

.lib 'C:\mdsy\rf018.l' TT
.END