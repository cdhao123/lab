
.PARAM VG = 1 VDD = 0.5 VDS = 5
M1 VIN VDD 0 0 N_1u L = 0.5U W = 1U
.INCLUDE 'C:\sdsy\model1\rf018.l'
VDD VDD 0 VDD
VIN VIN 0 VDS

.DC VIN 0 5 0.001

.PRINT i(M1) v(VIN)

.OPTION LIST NODE BRIEF=1 
.OPTION POST=3

.ALTER
.PARAM VDD = 1
.ALTER
.PARAM VDD = 1.5
.ALTER
.PARAM VDD = 2
.ALTER
.PARAM VDD = 2.5

.END