
.PARAM CLOAD = 0
M0 Z CLK 0 0 N_50n L = 50N W = 500N
M1 X A Z 0 N_50n L = 50N W = 500N
M2 Y B X 0 N_50n L = 50N W = 500N
M3 Y CLK VDD VDD P_50n L = 50N W = 250N
CL Y 0 2F

VCLK CLK 0 PULSE 0 1 4.995N 0.01N 0.01N 5N 10N
VDD VDD 0 1
VA A 0 PWL 0N 0 25N 0 14.99N 0 15N 1 19.99N 1 20N 0
VB B 0 PWL 0 0 5.99N 0 6N 1 12.99N 1 13N 0 14.99N 0 15N 1 19.99N 1 20N 0

.INCLUDE '..\model1\rf018.l'
* .DC VIN 0 1 0.001
.TRAN 0.001N 25N START = 0

.measure tran thl when V(Y) = 0.5 fall = 1
.measure tran tlh when V(Y) = 0.5 rise = 1

.OPTION LIST NODE BRIEF=1 
.OPTION POST=3

.END