
.PARAM VG = 1 VDD = 2.5 VDS = 5 LEN = 0.45U WID = 0.9U
M1 VIN VDD 0 0 N_1u L = LEN W = WID
.INCLUDE 'C:\sdsy\model1\rf018.l'
VDD VDD 0 VDD
VIN VIN 0 VDS

.DC VIN 0 5 0.001

.PRINT i(M1) v(VIN)

.OPTION LIST NODE BRIEF=1 
.OPTION POST=3

.ALTER
.PARAM LEN = 0.5U WID = 1U
.ALTER
.PARAM LEN = 0.55U WID = 1.1U
.ALTER
.PARAM LEN = 0.6U WID = 1.2U

.END