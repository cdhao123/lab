
.PARAM VDD = 1.8 WP = 5U
M1 VIN VIN VDD VDD PCH L = 0.18U W = WP
VDD VDD 0 VDD
VIN VIN 0 1

* .DC VIN 0 1.8 0.001
.DC WP 5U 10U 0.01U

.PRINT GM = par('LX7(M1)') IDS = par('LX4(M1)')

.OPTION LIST NODE BRIEF=1 
.OPTION POST=3

.lib 'C:\mdsy\rf018.l' TT
.END