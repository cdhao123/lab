
M0 VM0D VINB 0 0 N_50n L = 50N W = 0.5U
M1 VOUT VINA VM0D 0 N_50n L = 50N W = 0.5U
M2 VOUT VINA VDD VDD P_50n L = 50N W = 1U
M3 VOUT VINB VDD VDD P_50n L = 50N W = 1U

M4 VM4D VDD 0 0 N_50n L = 50N W = 0.5U
M5 VOUT2 VOUT VM4D 0 N_50n L = 50N W = 0.5U
M6 VOUT2 VOUT VDD VDD P_50n L = 50N W = 1U
M7 VOUT2 VDD VDD VDD P_50n L = 50N W = 1U

V1 VINA 0 1
V2 VINB 0 PULSE 0 1 10N 0.01N 0.01N 20N 40N

VDD VDD 0 1
.INCLUDE 'C:\sdsy\model1\rf018.l'
* .DC VINB 0 1 0.001
* .DC VINA 0 1 0.001
.TRAN 0.01N 40N START = 0
.measure tran thl when V(VOUT) = 0.5 fall = 1
.measure tran tlh when V(VOUT) = 0.5 rise = 1

.OPTION LIST NODE BRIEF=1 
.OPTION POST=3

.ALTER
V1 VINA 0 PULSE 0 1 10N 0.01N 0.01N 20N 40N
V2 VINB 0 1

.END