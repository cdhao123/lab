
.PARAM VDD = 1 R1 = 5000 VGS = 1 WP = 0.5U
M1 VOUT VIN 0 0 N_50n L = 0.05U W = 1U
M2 VOUT 0 VDD VDD P_50n L = 0.05U W = WP

.INCLUDE 'C:\sdsy\model1\rf018.l'

VDD VDD 0 VDD
VIN VIN 0 VGS

.DC VIN 0 1 0.001

.PRINT v(VIN) v(VOUT)

.OPTION LIST NODE BRIEF=1 
.OPTION POST=3

.ALTER
.PARAM WP = 1U

.END