* .PARAM VDD = 1 VGS = 1 LN = 0.05U LP = 0.05U WN = 1U WP = 0.5U
* M1 VOUT VIN 0 0 N_50n L = LN W = WN
* M2 VOUT VIN VDD VDD P_50n L = LP W = WP
* C1 
.PARAM VDD = 1.8
M1 VM1D VIN 0 0 NCH L = 0.25U W = 8U
M2 VM2D VIN VDD VDD PCH L = 0.25U W = 20U
V1 VM1D 0 0.2
V2 VM2D 0 1.6
VIN VIN 0 1.8

VDD VDD 0 VDD
.DC VIN 0 1.8 0.001

.PRINT i(VM1D) i(VM2D)
.PRINT M1_VTH = par('lv9(M1)')
.PRINT M2_VTH = par('lv9(M2)')


.OPTION LIST NODE BRIEF=1 
.OPTION POST=3

.lib 'C:\mdsy\rf018.l' TT
.END