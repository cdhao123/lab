
* .PARAM VDD = 1 VGS = 1 LN = 0.05U LP = 0.05U WN = 1U WP = 0.5U
* M1 VOUT VIN 0 0 N_50n L = LN W = WN
* M2 VOUT VIN VDD VDD P_50n L = LP W = WP
* C1 
.PARAM VDD = 1.8 NFACTOR = 1 PFACTOR = 1 VBIAS = 1.1517
I1 VDD VM2D 130U
* current mirror
M2 VM2D VM2D 0 0 NCH L = 1U W = 32U
M4 VB2 VM2D 0 0 NCH L = 1U W = 32U
M8 VB3 VM2D 0 0 NCH L = 1U W = 32U
* NMOS
M12 VB1 VB1 0 0 NCH L = NFACTOR*0.25U W = NFACTOR*1.6U
M15 VM15D VB4 0 0 NCH L = NFACTOR*0.25U W = NFACTOR*8U
M16 VB4 VB1 VM15D 0 NCH L = NFACTOR*0.25U W = NFACTOR*8U
M5 VM5D VB4 0 0 NCH L = NFACTOR*0.25U W = NFACTOR*16U
M3 VOUT VB1 VM5D 0 NCH L = NFACTOR*0.25U W = NFACTOR*8U
*PMOS
M6 VB2 VB2 VDD VDD PCH L = PFACTOR*0.25U W = PFACTOR*4U
M10 VB3 VB2 VM10S VDD PCH L = PFACTOR*0.25U W = PFACTOR*20U
M11 VM10S VB3 VDD VDD PCH L = PFACTOR*0.25U W = PFACTOR*20U
M13 VB1 VB2 VM13S VDD PCH L = PFACTOR*0.25U W = PFACTOR*20U
M14 VM13S VB3 VDD VDD PCH L = PFACTOR*0.25U W = PFACTOR*20U
M17 VB4 VB2 VM17S VDD PCH L = PFACTOR*0.25U W = PFACTOR*20U
M18 VM17S VB3 VDD VDD PCH L = PFACTOR*0.25U W = PFACTOR*20U
M7 VOUT VB2 VM7S VDD PCH L = PFACTOR*0.25U W = PFACTOR*20U
M9 VM7S VB3 VDD VDD PCH L = PFACTOR*0.25U W = PFACTOR*20U
M1 VM5D VIN VDD VDD PCH L = PFACTOR*0.18U W = PFACTOR*15U
C1 VOUT 0 5.0e-12


VDD VDD 0 VDD
* VIN VIN 0 PULSE (0 1 5NS 0.01NS 0.01NS 5NS)
VIN VIN 0 VBIAS AC = 1
* VOUTSIN VOUT 0 SIN VBIAS 1 10
* VOUT VOUT 0 VBIAS AC = 1


* .DC VIN 0 1.8 0.0001
.AC DEC 10 1 1G
* .DC VBIAS 0 1.8 0.001
* .TRAN 0.001NS 25NS START = 0S STOP = 25NS
* .measure tran tdlay1f trig V(VOUT) val=0.5 td=5n rise=1 targ V(VOUT) val=1 fall=1
* .measure tran thl when V(VOUT) = 0.5 fall = 1
* .measure tran tlh when V(VOUT) = 0.5 rise = 1
* .PRINT v(VIN) v(VOUT)


.lib 'C:\mdsy\rf018.l' TT

.OPTION LIST NODE BRIEF=1 
.OPTION POST=3

.ALTER
.PARAM NFACTOR = 2 VBIAS = 1.154
.ALTER
.PARAM NFACTOR = 4 VBIAS = 1.154
.ALTER
.PARAM NFACTOR = 8 VBIAS = 1.1548
.ALTER
.PARAM NFACTOR = 16 VBIAS = 1.1548
.ALTER
.PARAM NFACTOR = 16 PFACTOR = 2 VBIAS = 1.1415
.ALTER
.PARAM NFACTOR = 16 PFACTOR = 4 VBIAS = 1.1351
.ALTER
.PARAM NFACTOR = 16 PFACTOR = 8 VBIAS = 1.1373

.END