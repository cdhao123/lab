
.PARAM VG = 1 VDD = 0.7 VDS = 5
M1 0 VDD VIN 0 P_50n L = 0.05U W = 0.1U
.INCLUDE 'C:\sdsy\model1\rf018.l'
VDD VDD 0 VDD
VIN VIN 0 VDS

.DC VIN 0 1 0.001

.PRINT i(M1) v(VIN)

.OPTION LIST NODE BRIEF=1 
.OPTION POST=3

.ALTER
.PARAM VDD = 0.8
.ALTER
.PARAM VDD = 0.9
.ALTER
.PARAM VDD = 0.95
.ALTER
.PARAM VDD = 1

.END