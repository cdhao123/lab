
* .PARAM VDD = 1 VGS = 1 LN = 0.05U LP = 0.05U WN = 1U WP = 0.5U
* M1 VOUT VIN 0 0 N_50n L = LN W = WN
* M2 VOUT VIN VDD VDD P_50n L = LP W = WP
* C1 
.PARAM VDD = 1 LN = 0.05U LP = 0.05U WN = 0.05U WP = 0.075U A = 3.51
M1 VOUT1 VIN 0 0 N_50n L = LN W = WN
M2 VOUT1 VIN VDD VDD P_50n L = LP W = WP
M3 VOUT2 VOUT1 0 0 N_50n L = 0.05U W = A*WN
M4 VOUT2 VOUT1 VDD VDD P_50n L = 0.075U W = A*WP
M5 VOUT3 VOUT2 0 0 N_50n L = 0.05U W = A*A*WN
M6 VOUT3 VOUT2 VDD VDD P_50n L = 0.075U W = A*A*WP
M7 VOUT4 VOUT3 0 0 N_50n L = 0.05U W = A*A*A*WN
M8 VOUT4 VOUT3 VDD VDD P_50n L = 0.075U W = A*A*A*WP
* M9  VOUT5 VOUT4 0 0 N_50n L = 0.05U W = A*A*A*A*WN
* M10 VOUT5 VOUT4 VDD VDD P_50n L = 0.075U W = A*A*A*A*WP
* M11 VOUT6 VOUT5 0 0 N_50n L = 0.05U W = A*A*A*A*A*WN
* M12 VOUT6 VOUT5 VDD VDD P_50n L = 0.075U W = A*A*A*A*A*WP
* M13 VOUT7 VOUT6 0 0 N_50n L = 0.05U W = A*A*A*A*A*A*WN
* M14 VOUT7 VOUT6 VDD VDD P_50n L = 0.075U W = A*A*A*A*A*A*WP
C1 VOUT4 0 5.0e-12
.INCLUDE 'C:\sdsy\model1\rf018.l'

VDD VDD 0 VDD
VIN VIN 0 PULSE (0 1 5NS 0.01NS 0.01NS 40NS)

.TRAN 0.001NS 60NS START = 0S STOP = 60NS
* .measure tran tdlay1f trig V(VOUT) val=0.5 td=5n rise=1 targ V(VOUT) val=1 fall=1
.measure tran thl when V(VOUT4) = 0.5 fall = 1
.measure tran tlh when V(VOUT4) = 0.5 rise = 1
.PRINT v(VIN) v(VOUT4)



.OPTION LIST NODE BRIEF=1 
.OPTION POST=3

.END